library ads;
use ads.ads_fixed.all;
use ads.ads_complex_pkg.all;

package seed_table is
	type seed_rom_type is array (natural range<>) of ads_complex;
	constant seed_rom: seed_rom_type := (
			( re => to_ads_sfixed( 0.75000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed( 0.74992), im => to_ads_sfixed( 0.01122) ),
			( re => to_ads_sfixed( 0.74966), im => to_ads_sfixed( 0.02244) ),
			( re => to_ads_sfixed( 0.74924), im => to_ads_sfixed( 0.03365) ),
			( re => to_ads_sfixed( 0.74866), im => to_ads_sfixed( 0.04485) ),
			( re => to_ads_sfixed( 0.74790), im => to_ads_sfixed( 0.05605) ),
			( re => to_ads_sfixed( 0.74698), im => to_ads_sfixed( 0.06723) ),
			( re => to_ads_sfixed( 0.74589), im => to_ads_sfixed( 0.07840) ),
			( re => to_ads_sfixed( 0.74464), im => to_ads_sfixed( 0.08955) ),
			( re => to_ads_sfixed( 0.74321), im => to_ads_sfixed( 0.10067) ),
			( re => to_ads_sfixed( 0.74162), im => to_ads_sfixed( 0.11178) ),
			( re => to_ads_sfixed( 0.73987), im => to_ads_sfixed( 0.12286) ),
			( re => to_ads_sfixed( 0.73795), im => to_ads_sfixed( 0.13392) ),
			( re => to_ads_sfixed( 0.73586), im => to_ads_sfixed( 0.14494) ),
			( re => to_ads_sfixed( 0.73361), im => to_ads_sfixed( 0.15593) ),
			( re => to_ads_sfixed( 0.73120), im => to_ads_sfixed( 0.16689) ),
			( re => to_ads_sfixed( 0.72862), im => to_ads_sfixed( 0.17781) ),
			( re => to_ads_sfixed( 0.72588), im => to_ads_sfixed( 0.18869) ),
			( re => to_ads_sfixed( 0.72297), im => to_ads_sfixed( 0.19953) ),
			( re => to_ads_sfixed( 0.71991), im => to_ads_sfixed( 0.21032) ),
			( re => to_ads_sfixed( 0.71668), im => to_ads_sfixed( 0.22107) ),
			( re => to_ads_sfixed( 0.71329), im => to_ads_sfixed( 0.23176) ),
			( re => to_ads_sfixed( 0.70975), im => to_ads_sfixed( 0.24241) ),
			( re => to_ads_sfixed( 0.70604), im => to_ads_sfixed( 0.25300) ),
			( re => to_ads_sfixed( 0.70218), im => to_ads_sfixed( 0.26353) ),
			( re => to_ads_sfixed( 0.69816), im => to_ads_sfixed( 0.27401) ),
			( re => to_ads_sfixed( 0.69398), im => to_ads_sfixed( 0.28442) ),
			( re => to_ads_sfixed( 0.68965), im => to_ads_sfixed( 0.29477) ),
			( re => to_ads_sfixed( 0.68516), im => to_ads_sfixed( 0.30505) ),
			( re => to_ads_sfixed( 0.68052), im => to_ads_sfixed( 0.31527) ),
			( re => to_ads_sfixed( 0.67573), im => to_ads_sfixed( 0.32541) ),
			( re => to_ads_sfixed( 0.67078), im => to_ads_sfixed( 0.33548) ),
			( re => to_ads_sfixed( 0.66569), im => to_ads_sfixed( 0.34548) ),
			( re => to_ads_sfixed( 0.66045), im => to_ads_sfixed( 0.35540) ),
			( re => to_ads_sfixed( 0.65506), im => to_ads_sfixed( 0.36524) ),
			( re => to_ads_sfixed( 0.64952), im => to_ads_sfixed( 0.37500) ),
			( re => to_ads_sfixed( 0.64384), im => to_ads_sfixed( 0.38467) ),
			( re => to_ads_sfixed( 0.63801), im => to_ads_sfixed( 0.39426) ),
			( re => to_ads_sfixed( 0.63204), im => to_ads_sfixed( 0.40376) ),
			( re => to_ads_sfixed( 0.62593), im => to_ads_sfixed( 0.41317) ),
			( re => to_ads_sfixed( 0.61968), im => to_ads_sfixed( 0.42249) ),
			( re => to_ads_sfixed( 0.61329), im => to_ads_sfixed( 0.43171) ),
			( re => to_ads_sfixed( 0.60676), im => to_ads_sfixed( 0.44084) ),
			( re => to_ads_sfixed( 0.60010), im => to_ads_sfixed( 0.44987) ),
			( re => to_ads_sfixed( 0.59330), im => to_ads_sfixed( 0.45879) ),
			( re => to_ads_sfixed( 0.58637), im => to_ads_sfixed( 0.46762) ),
			( re => to_ads_sfixed( 0.57931), im => to_ads_sfixed( 0.47634) ),
			( re => to_ads_sfixed( 0.57212), im => to_ads_sfixed( 0.48495) ),
			( re => to_ads_sfixed( 0.56480), im => to_ads_sfixed( 0.49345) ),
			( re => to_ads_sfixed( 0.55736), im => to_ads_sfixed( 0.50185) ),
			( re => to_ads_sfixed( 0.54979), im => to_ads_sfixed( 0.51013) ),
			( re => to_ads_sfixed( 0.54210), im => to_ads_sfixed( 0.51830) ),
			( re => to_ads_sfixed( 0.53428), im => to_ads_sfixed( 0.52635) ),
			( re => to_ads_sfixed( 0.52635), im => to_ads_sfixed( 0.53428) ),
			( re => to_ads_sfixed( 0.51830), im => to_ads_sfixed( 0.54210) ),
			( re => to_ads_sfixed( 0.51013), im => to_ads_sfixed( 0.54979) ),
			( re => to_ads_sfixed( 0.50185), im => to_ads_sfixed( 0.55736) ),
			( re => to_ads_sfixed( 0.49345), im => to_ads_sfixed( 0.56480) ),
			( re => to_ads_sfixed( 0.48495), im => to_ads_sfixed( 0.57212) ),
			( re => to_ads_sfixed( 0.47634), im => to_ads_sfixed( 0.57931) ),
			( re => to_ads_sfixed( 0.46762), im => to_ads_sfixed( 0.58637) ),
			( re => to_ads_sfixed( 0.45879), im => to_ads_sfixed( 0.59330) ),
			( re => to_ads_sfixed( 0.44987), im => to_ads_sfixed( 0.60010) ),
			( re => to_ads_sfixed( 0.44084), im => to_ads_sfixed( 0.60676) ),
			( re => to_ads_sfixed( 0.43171), im => to_ads_sfixed( 0.61329) ),
			( re => to_ads_sfixed( 0.42249), im => to_ads_sfixed( 0.61968) ),
			( re => to_ads_sfixed( 0.41317), im => to_ads_sfixed( 0.62593) ),
			( re => to_ads_sfixed( 0.40376), im => to_ads_sfixed( 0.63204) ),
			( re => to_ads_sfixed( 0.39426), im => to_ads_sfixed( 0.63801) ),
			( re => to_ads_sfixed( 0.38467), im => to_ads_sfixed( 0.64384) ),
			( re => to_ads_sfixed( 0.37500), im => to_ads_sfixed( 0.64952) ),
			( re => to_ads_sfixed( 0.36524), im => to_ads_sfixed( 0.65506) ),
			( re => to_ads_sfixed( 0.35540), im => to_ads_sfixed( 0.66045) ),
			( re => to_ads_sfixed( 0.34548), im => to_ads_sfixed( 0.66569) ),
			( re => to_ads_sfixed( 0.33548), im => to_ads_sfixed( 0.67078) ),
			( re => to_ads_sfixed( 0.32541), im => to_ads_sfixed( 0.67573) ),
			( re => to_ads_sfixed( 0.31527), im => to_ads_sfixed( 0.68052) ),
			( re => to_ads_sfixed( 0.30505), im => to_ads_sfixed( 0.68516) ),
			( re => to_ads_sfixed( 0.29477), im => to_ads_sfixed( 0.68965) ),
			( re => to_ads_sfixed( 0.28442), im => to_ads_sfixed( 0.69398) ),
			( re => to_ads_sfixed( 0.27401), im => to_ads_sfixed( 0.69816) ),
			( re => to_ads_sfixed( 0.26353), im => to_ads_sfixed( 0.70218) ),
			( re => to_ads_sfixed( 0.25300), im => to_ads_sfixed( 0.70604) ),
			( re => to_ads_sfixed( 0.24241), im => to_ads_sfixed( 0.70975) ),
			( re => to_ads_sfixed( 0.23176), im => to_ads_sfixed( 0.71329) ),
			( re => to_ads_sfixed( 0.22107), im => to_ads_sfixed( 0.71668) ),
			( re => to_ads_sfixed( 0.21032), im => to_ads_sfixed( 0.71991) ),
			( re => to_ads_sfixed( 0.19953), im => to_ads_sfixed( 0.72297) ),
			( re => to_ads_sfixed( 0.18869), im => to_ads_sfixed( 0.72588) ),
			( re => to_ads_sfixed( 0.17781), im => to_ads_sfixed( 0.72862) ),
			( re => to_ads_sfixed( 0.16689), im => to_ads_sfixed( 0.73120) ),
			( re => to_ads_sfixed( 0.15593), im => to_ads_sfixed( 0.73361) ),
			( re => to_ads_sfixed( 0.14494), im => to_ads_sfixed( 0.73586) ),
			( re => to_ads_sfixed( 0.13392), im => to_ads_sfixed( 0.73795) ),
			( re => to_ads_sfixed( 0.12286), im => to_ads_sfixed( 0.73987) ),
			( re => to_ads_sfixed( 0.11178), im => to_ads_sfixed( 0.74162) ),
			( re => to_ads_sfixed( 0.10067), im => to_ads_sfixed( 0.74321) ),
			( re => to_ads_sfixed( 0.08955), im => to_ads_sfixed( 0.74464) ),
			( re => to_ads_sfixed( 0.07840), im => to_ads_sfixed( 0.74589) ),
			( re => to_ads_sfixed( 0.06723), im => to_ads_sfixed( 0.74698) ),
			( re => to_ads_sfixed( 0.05605), im => to_ads_sfixed( 0.74790) ),
			( re => to_ads_sfixed( 0.04485), im => to_ads_sfixed( 0.74866) ),
			( re => to_ads_sfixed( 0.03365), im => to_ads_sfixed( 0.74924) ),
			( re => to_ads_sfixed( 0.02244), im => to_ads_sfixed( 0.74966) ),
			( re => to_ads_sfixed( 0.01122), im => to_ads_sfixed( 0.74992) ),
			( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed( 0.75000) ),
			( re => to_ads_sfixed(-0.01122), im => to_ads_sfixed( 0.74992) ),
			( re => to_ads_sfixed(-0.02244), im => to_ads_sfixed( 0.74966) ),
			( re => to_ads_sfixed(-0.03365), im => to_ads_sfixed( 0.74924) ),
			( re => to_ads_sfixed(-0.04485), im => to_ads_sfixed( 0.74866) ),
			( re => to_ads_sfixed(-0.05605), im => to_ads_sfixed( 0.74790) ),
			( re => to_ads_sfixed(-0.06723), im => to_ads_sfixed( 0.74698) ),
			( re => to_ads_sfixed(-0.07840), im => to_ads_sfixed( 0.74589) ),
			( re => to_ads_sfixed(-0.08955), im => to_ads_sfixed( 0.74464) ),
			( re => to_ads_sfixed(-0.10067), im => to_ads_sfixed( 0.74321) ),
			( re => to_ads_sfixed(-0.11178), im => to_ads_sfixed( 0.74162) ),
			( re => to_ads_sfixed(-0.12286), im => to_ads_sfixed( 0.73987) ),
			( re => to_ads_sfixed(-0.13392), im => to_ads_sfixed( 0.73795) ),
			( re => to_ads_sfixed(-0.14494), im => to_ads_sfixed( 0.73586) ),
			( re => to_ads_sfixed(-0.15593), im => to_ads_sfixed( 0.73361) ),
			( re => to_ads_sfixed(-0.16689), im => to_ads_sfixed( 0.73120) ),
			( re => to_ads_sfixed(-0.17781), im => to_ads_sfixed( 0.72862) ),
			( re => to_ads_sfixed(-0.18869), im => to_ads_sfixed( 0.72588) ),
			( re => to_ads_sfixed(-0.19953), im => to_ads_sfixed( 0.72297) ),
			( re => to_ads_sfixed(-0.21032), im => to_ads_sfixed( 0.71991) ),
			( re => to_ads_sfixed(-0.22107), im => to_ads_sfixed( 0.71668) ),
			( re => to_ads_sfixed(-0.23176), im => to_ads_sfixed( 0.71329) ),
			( re => to_ads_sfixed(-0.24241), im => to_ads_sfixed( 0.70975) ),
			( re => to_ads_sfixed(-0.25300), im => to_ads_sfixed( 0.70604) ),
			( re => to_ads_sfixed(-0.26353), im => to_ads_sfixed( 0.70218) ),
			( re => to_ads_sfixed(-0.27401), im => to_ads_sfixed( 0.69816) ),
			( re => to_ads_sfixed(-0.28442), im => to_ads_sfixed( 0.69398) ),
			( re => to_ads_sfixed(-0.29477), im => to_ads_sfixed( 0.68965) ),
			( re => to_ads_sfixed(-0.30505), im => to_ads_sfixed( 0.68516) ),
			( re => to_ads_sfixed(-0.31527), im => to_ads_sfixed( 0.68052) ),
			( re => to_ads_sfixed(-0.32541), im => to_ads_sfixed( 0.67573) ),
			( re => to_ads_sfixed(-0.33548), im => to_ads_sfixed( 0.67078) ),
			( re => to_ads_sfixed(-0.34548), im => to_ads_sfixed( 0.66569) ),
			( re => to_ads_sfixed(-0.35540), im => to_ads_sfixed( 0.66045) ),
			( re => to_ads_sfixed(-0.36524), im => to_ads_sfixed( 0.65506) ),
			( re => to_ads_sfixed(-0.37500), im => to_ads_sfixed( 0.64952) ),
			( re => to_ads_sfixed(-0.38467), im => to_ads_sfixed( 0.64384) ),
			( re => to_ads_sfixed(-0.39426), im => to_ads_sfixed( 0.63801) ),
			( re => to_ads_sfixed(-0.40376), im => to_ads_sfixed( 0.63204) ),
			( re => to_ads_sfixed(-0.41317), im => to_ads_sfixed( 0.62593) ),
			( re => to_ads_sfixed(-0.42249), im => to_ads_sfixed( 0.61968) ),
			( re => to_ads_sfixed(-0.43171), im => to_ads_sfixed( 0.61329) ),
			( re => to_ads_sfixed(-0.44084), im => to_ads_sfixed( 0.60676) ),
			( re => to_ads_sfixed(-0.44987), im => to_ads_sfixed( 0.60010) ),
			( re => to_ads_sfixed(-0.45879), im => to_ads_sfixed( 0.59330) ),
			( re => to_ads_sfixed(-0.46762), im => to_ads_sfixed( 0.58637) ),
			( re => to_ads_sfixed(-0.47634), im => to_ads_sfixed( 0.57931) ),
			( re => to_ads_sfixed(-0.48495), im => to_ads_sfixed( 0.57212) ),
			( re => to_ads_sfixed(-0.49345), im => to_ads_sfixed( 0.56480) ),
			( re => to_ads_sfixed(-0.50185), im => to_ads_sfixed( 0.55736) ),
			( re => to_ads_sfixed(-0.51013), im => to_ads_sfixed( 0.54979) ),
			( re => to_ads_sfixed(-0.51830), im => to_ads_sfixed( 0.54210) ),
			( re => to_ads_sfixed(-0.52635), im => to_ads_sfixed( 0.53428) ),
			( re => to_ads_sfixed(-0.53428), im => to_ads_sfixed( 0.52635) ),
			( re => to_ads_sfixed(-0.54210), im => to_ads_sfixed( 0.51830) ),
			( re => to_ads_sfixed(-0.54979), im => to_ads_sfixed( 0.51013) ),
			( re => to_ads_sfixed(-0.55736), im => to_ads_sfixed( 0.50185) ),
			( re => to_ads_sfixed(-0.56480), im => to_ads_sfixed( 0.49345) ),
			( re => to_ads_sfixed(-0.57212), im => to_ads_sfixed( 0.48495) ),
			( re => to_ads_sfixed(-0.57931), im => to_ads_sfixed( 0.47634) ),
			( re => to_ads_sfixed(-0.58637), im => to_ads_sfixed( 0.46762) ),
			( re => to_ads_sfixed(-0.59330), im => to_ads_sfixed( 0.45879) ),
			( re => to_ads_sfixed(-0.60010), im => to_ads_sfixed( 0.44987) ),
			( re => to_ads_sfixed(-0.60676), im => to_ads_sfixed( 0.44084) ),
			( re => to_ads_sfixed(-0.61329), im => to_ads_sfixed( 0.43171) ),
			( re => to_ads_sfixed(-0.61968), im => to_ads_sfixed( 0.42249) ),
			( re => to_ads_sfixed(-0.62593), im => to_ads_sfixed( 0.41317) ),
			( re => to_ads_sfixed(-0.63204), im => to_ads_sfixed( 0.40376) ),
			( re => to_ads_sfixed(-0.63801), im => to_ads_sfixed( 0.39426) ),
			( re => to_ads_sfixed(-0.64384), im => to_ads_sfixed( 0.38467) ),
			( re => to_ads_sfixed(-0.64952), im => to_ads_sfixed( 0.37500) ),
			( re => to_ads_sfixed(-0.65506), im => to_ads_sfixed( 0.36524) ),
			( re => to_ads_sfixed(-0.66045), im => to_ads_sfixed( 0.35540) ),
			( re => to_ads_sfixed(-0.66569), im => to_ads_sfixed( 0.34548) ),
			( re => to_ads_sfixed(-0.67078), im => to_ads_sfixed( 0.33548) ),
			( re => to_ads_sfixed(-0.67573), im => to_ads_sfixed( 0.32541) ),
			( re => to_ads_sfixed(-0.68052), im => to_ads_sfixed( 0.31527) ),
			( re => to_ads_sfixed(-0.68516), im => to_ads_sfixed( 0.30505) ),
			( re => to_ads_sfixed(-0.68965), im => to_ads_sfixed( 0.29477) ),
			( re => to_ads_sfixed(-0.69398), im => to_ads_sfixed( 0.28442) ),
			( re => to_ads_sfixed(-0.69816), im => to_ads_sfixed( 0.27401) ),
			( re => to_ads_sfixed(-0.70218), im => to_ads_sfixed( 0.26353) ),
			( re => to_ads_sfixed(-0.70604), im => to_ads_sfixed( 0.25300) ),
			( re => to_ads_sfixed(-0.70975), im => to_ads_sfixed( 0.24241) ),
			( re => to_ads_sfixed(-0.71329), im => to_ads_sfixed( 0.23176) ),
			( re => to_ads_sfixed(-0.71668), im => to_ads_sfixed( 0.22107) ),
			( re => to_ads_sfixed(-0.71991), im => to_ads_sfixed( 0.21032) ),
			( re => to_ads_sfixed(-0.72297), im => to_ads_sfixed( 0.19953) ),
			( re => to_ads_sfixed(-0.72588), im => to_ads_sfixed( 0.18869) ),
			( re => to_ads_sfixed(-0.72862), im => to_ads_sfixed( 0.17781) ),
			( re => to_ads_sfixed(-0.73120), im => to_ads_sfixed( 0.16689) ),
			( re => to_ads_sfixed(-0.73361), im => to_ads_sfixed( 0.15593) ),
			( re => to_ads_sfixed(-0.73586), im => to_ads_sfixed( 0.14494) ),
			( re => to_ads_sfixed(-0.73795), im => to_ads_sfixed( 0.13392) ),
			( re => to_ads_sfixed(-0.73987), im => to_ads_sfixed( 0.12286) ),
			( re => to_ads_sfixed(-0.74162), im => to_ads_sfixed( 0.11178) ),
			( re => to_ads_sfixed(-0.74321), im => to_ads_sfixed( 0.10067) ),
			( re => to_ads_sfixed(-0.74464), im => to_ads_sfixed( 0.08955) ),
			( re => to_ads_sfixed(-0.74589), im => to_ads_sfixed( 0.07840) ),
			( re => to_ads_sfixed(-0.74698), im => to_ads_sfixed( 0.06723) ),
			( re => to_ads_sfixed(-0.74790), im => to_ads_sfixed( 0.05605) ),
			( re => to_ads_sfixed(-0.74866), im => to_ads_sfixed( 0.04485) ),
			( re => to_ads_sfixed(-0.74924), im => to_ads_sfixed( 0.03365) ),
			( re => to_ads_sfixed(-0.74966), im => to_ads_sfixed( 0.02244) ),
			( re => to_ads_sfixed(-0.74992), im => to_ads_sfixed( 0.01122) ),
			( re => to_ads_sfixed(-0.75000), im => to_ads_sfixed(-0.00000) ),
			( re => to_ads_sfixed(-0.74992), im => to_ads_sfixed(-0.01122) ),
			( re => to_ads_sfixed(-0.74966), im => to_ads_sfixed(-0.02244) ),
			( re => to_ads_sfixed(-0.74924), im => to_ads_sfixed(-0.03365) ),
			( re => to_ads_sfixed(-0.74866), im => to_ads_sfixed(-0.04485) ),
			( re => to_ads_sfixed(-0.74790), im => to_ads_sfixed(-0.05605) ),
			( re => to_ads_sfixed(-0.74698), im => to_ads_sfixed(-0.06723) ),
			( re => to_ads_sfixed(-0.74589), im => to_ads_sfixed(-0.07840) ),
			( re => to_ads_sfixed(-0.74464), im => to_ads_sfixed(-0.08955) ),
			( re => to_ads_sfixed(-0.74321), im => to_ads_sfixed(-0.10067) ),
			( re => to_ads_sfixed(-0.74162), im => to_ads_sfixed(-0.11178) ),
			( re => to_ads_sfixed(-0.73987), im => to_ads_sfixed(-0.12286) ),
			( re => to_ads_sfixed(-0.73795), im => to_ads_sfixed(-0.13392) ),
			( re => to_ads_sfixed(-0.73586), im => to_ads_sfixed(-0.14494) ),
			( re => to_ads_sfixed(-0.73361), im => to_ads_sfixed(-0.15593) ),
			( re => to_ads_sfixed(-0.73120), im => to_ads_sfixed(-0.16689) ),
			( re => to_ads_sfixed(-0.72862), im => to_ads_sfixed(-0.17781) ),
			( re => to_ads_sfixed(-0.72588), im => to_ads_sfixed(-0.18869) ),
			( re => to_ads_sfixed(-0.72297), im => to_ads_sfixed(-0.19953) ),
			( re => to_ads_sfixed(-0.71991), im => to_ads_sfixed(-0.21032) ),
			( re => to_ads_sfixed(-0.71668), im => to_ads_sfixed(-0.22107) ),
			( re => to_ads_sfixed(-0.71329), im => to_ads_sfixed(-0.23176) ),
			( re => to_ads_sfixed(-0.70975), im => to_ads_sfixed(-0.24241) ),
			( re => to_ads_sfixed(-0.70604), im => to_ads_sfixed(-0.25300) ),
			( re => to_ads_sfixed(-0.70218), im => to_ads_sfixed(-0.26353) ),
			( re => to_ads_sfixed(-0.69816), im => to_ads_sfixed(-0.27401) ),
			( re => to_ads_sfixed(-0.69398), im => to_ads_sfixed(-0.28442) ),
			( re => to_ads_sfixed(-0.68965), im => to_ads_sfixed(-0.29477) ),
			( re => to_ads_sfixed(-0.68516), im => to_ads_sfixed(-0.30505) ),
			( re => to_ads_sfixed(-0.68052), im => to_ads_sfixed(-0.31527) ),
			( re => to_ads_sfixed(-0.67573), im => to_ads_sfixed(-0.32541) ),
			( re => to_ads_sfixed(-0.67078), im => to_ads_sfixed(-0.33548) ),
			( re => to_ads_sfixed(-0.66569), im => to_ads_sfixed(-0.34548) ),
			( re => to_ads_sfixed(-0.66045), im => to_ads_sfixed(-0.35540) ),
			( re => to_ads_sfixed(-0.65506), im => to_ads_sfixed(-0.36524) ),
			( re => to_ads_sfixed(-0.64952), im => to_ads_sfixed(-0.37500) ),
			( re => to_ads_sfixed(-0.64384), im => to_ads_sfixed(-0.38467) ),
			( re => to_ads_sfixed(-0.63801), im => to_ads_sfixed(-0.39426) ),
			( re => to_ads_sfixed(-0.63204), im => to_ads_sfixed(-0.40376) ),
			( re => to_ads_sfixed(-0.62593), im => to_ads_sfixed(-0.41317) ),
			( re => to_ads_sfixed(-0.61968), im => to_ads_sfixed(-0.42249) ),
			( re => to_ads_sfixed(-0.61329), im => to_ads_sfixed(-0.43171) ),
			( re => to_ads_sfixed(-0.60676), im => to_ads_sfixed(-0.44084) ),
			( re => to_ads_sfixed(-0.60010), im => to_ads_sfixed(-0.44987) ),
			( re => to_ads_sfixed(-0.59330), im => to_ads_sfixed(-0.45879) ),
			( re => to_ads_sfixed(-0.58637), im => to_ads_sfixed(-0.46762) ),
			( re => to_ads_sfixed(-0.57931), im => to_ads_sfixed(-0.47634) ),
			( re => to_ads_sfixed(-0.57212), im => to_ads_sfixed(-0.48495) ),
			( re => to_ads_sfixed(-0.56480), im => to_ads_sfixed(-0.49345) ),
			( re => to_ads_sfixed(-0.55736), im => to_ads_sfixed(-0.50185) ),
			( re => to_ads_sfixed(-0.54979), im => to_ads_sfixed(-0.51013) ),
			( re => to_ads_sfixed(-0.54210), im => to_ads_sfixed(-0.51830) ),
			( re => to_ads_sfixed(-0.53428), im => to_ads_sfixed(-0.52635) ),
			( re => to_ads_sfixed(-0.52635), im => to_ads_sfixed(-0.53428) ),
			( re => to_ads_sfixed(-0.51830), im => to_ads_sfixed(-0.54210) ),
			( re => to_ads_sfixed(-0.51013), im => to_ads_sfixed(-0.54979) ),
			( re => to_ads_sfixed(-0.50185), im => to_ads_sfixed(-0.55736) ),
			( re => to_ads_sfixed(-0.49345), im => to_ads_sfixed(-0.56480) ),
			( re => to_ads_sfixed(-0.48495), im => to_ads_sfixed(-0.57212) ),
			( re => to_ads_sfixed(-0.47634), im => to_ads_sfixed(-0.57931) ),
			( re => to_ads_sfixed(-0.46762), im => to_ads_sfixed(-0.58637) ),
			( re => to_ads_sfixed(-0.45879), im => to_ads_sfixed(-0.59330) ),
			( re => to_ads_sfixed(-0.44987), im => to_ads_sfixed(-0.60010) ),
			( re => to_ads_sfixed(-0.44084), im => to_ads_sfixed(-0.60676) ),
			( re => to_ads_sfixed(-0.43171), im => to_ads_sfixed(-0.61329) ),
			( re => to_ads_sfixed(-0.42249), im => to_ads_sfixed(-0.61968) ),
			( re => to_ads_sfixed(-0.41317), im => to_ads_sfixed(-0.62593) ),
			( re => to_ads_sfixed(-0.40376), im => to_ads_sfixed(-0.63204) ),
			( re => to_ads_sfixed(-0.39426), im => to_ads_sfixed(-0.63801) ),
			( re => to_ads_sfixed(-0.38467), im => to_ads_sfixed(-0.64384) ),
			( re => to_ads_sfixed(-0.37500), im => to_ads_sfixed(-0.64952) ),
			( re => to_ads_sfixed(-0.36524), im => to_ads_sfixed(-0.65506) ),
			( re => to_ads_sfixed(-0.35540), im => to_ads_sfixed(-0.66045) ),
			( re => to_ads_sfixed(-0.34548), im => to_ads_sfixed(-0.66569) ),
			( re => to_ads_sfixed(-0.33548), im => to_ads_sfixed(-0.67078) ),
			( re => to_ads_sfixed(-0.32541), im => to_ads_sfixed(-0.67573) ),
			( re => to_ads_sfixed(-0.31527), im => to_ads_sfixed(-0.68052) ),
			( re => to_ads_sfixed(-0.30505), im => to_ads_sfixed(-0.68516) ),
			( re => to_ads_sfixed(-0.29477), im => to_ads_sfixed(-0.68965) ),
			( re => to_ads_sfixed(-0.28442), im => to_ads_sfixed(-0.69398) ),
			( re => to_ads_sfixed(-0.27401), im => to_ads_sfixed(-0.69816) ),
			( re => to_ads_sfixed(-0.26353), im => to_ads_sfixed(-0.70218) ),
			( re => to_ads_sfixed(-0.25300), im => to_ads_sfixed(-0.70604) ),
			( re => to_ads_sfixed(-0.24241), im => to_ads_sfixed(-0.70975) ),
			( re => to_ads_sfixed(-0.23176), im => to_ads_sfixed(-0.71329) ),
			( re => to_ads_sfixed(-0.22107), im => to_ads_sfixed(-0.71668) ),
			( re => to_ads_sfixed(-0.21032), im => to_ads_sfixed(-0.71991) ),
			( re => to_ads_sfixed(-0.19953), im => to_ads_sfixed(-0.72297) ),
			( re => to_ads_sfixed(-0.18869), im => to_ads_sfixed(-0.72588) ),
			( re => to_ads_sfixed(-0.17781), im => to_ads_sfixed(-0.72862) ),
			( re => to_ads_sfixed(-0.16689), im => to_ads_sfixed(-0.73120) ),
			( re => to_ads_sfixed(-0.15593), im => to_ads_sfixed(-0.73361) ),
			( re => to_ads_sfixed(-0.14494), im => to_ads_sfixed(-0.73586) ),
			( re => to_ads_sfixed(-0.13392), im => to_ads_sfixed(-0.73795) ),
			( re => to_ads_sfixed(-0.12286), im => to_ads_sfixed(-0.73987) ),
			( re => to_ads_sfixed(-0.11178), im => to_ads_sfixed(-0.74162) ),
			( re => to_ads_sfixed(-0.10067), im => to_ads_sfixed(-0.74321) ),
			( re => to_ads_sfixed(-0.08955), im => to_ads_sfixed(-0.74464) ),
			( re => to_ads_sfixed(-0.07840), im => to_ads_sfixed(-0.74589) ),
			( re => to_ads_sfixed(-0.06723), im => to_ads_sfixed(-0.74698) ),
			( re => to_ads_sfixed(-0.05605), im => to_ads_sfixed(-0.74790) ),
			( re => to_ads_sfixed(-0.04485), im => to_ads_sfixed(-0.74866) ),
			( re => to_ads_sfixed(-0.03365), im => to_ads_sfixed(-0.74924) ),
			( re => to_ads_sfixed(-0.02244), im => to_ads_sfixed(-0.74966) ),
			( re => to_ads_sfixed(-0.01122), im => to_ads_sfixed(-0.74992) ),
			( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed(-0.75000) ),
			( re => to_ads_sfixed( 0.01122), im => to_ads_sfixed(-0.74992) ),
			( re => to_ads_sfixed( 0.02244), im => to_ads_sfixed(-0.74966) ),
			( re => to_ads_sfixed( 0.03365), im => to_ads_sfixed(-0.74924) ),
			( re => to_ads_sfixed( 0.04485), im => to_ads_sfixed(-0.74866) ),
			( re => to_ads_sfixed( 0.05605), im => to_ads_sfixed(-0.74790) ),
			( re => to_ads_sfixed( 0.06723), im => to_ads_sfixed(-0.74698) ),
			( re => to_ads_sfixed( 0.07840), im => to_ads_sfixed(-0.74589) ),
			( re => to_ads_sfixed( 0.08955), im => to_ads_sfixed(-0.74464) ),
			( re => to_ads_sfixed( 0.10067), im => to_ads_sfixed(-0.74321) ),
			( re => to_ads_sfixed( 0.11178), im => to_ads_sfixed(-0.74162) ),
			( re => to_ads_sfixed( 0.12286), im => to_ads_sfixed(-0.73987) ),
			( re => to_ads_sfixed( 0.13392), im => to_ads_sfixed(-0.73795) ),
			( re => to_ads_sfixed( 0.14494), im => to_ads_sfixed(-0.73586) ),
			( re => to_ads_sfixed( 0.15593), im => to_ads_sfixed(-0.73361) ),
			( re => to_ads_sfixed( 0.16689), im => to_ads_sfixed(-0.73120) ),
			( re => to_ads_sfixed( 0.17781), im => to_ads_sfixed(-0.72862) ),
			( re => to_ads_sfixed( 0.18869), im => to_ads_sfixed(-0.72588) ),
			( re => to_ads_sfixed( 0.19953), im => to_ads_sfixed(-0.72297) ),
			( re => to_ads_sfixed( 0.21032), im => to_ads_sfixed(-0.71991) ),
			( re => to_ads_sfixed( 0.22107), im => to_ads_sfixed(-0.71668) ),
			( re => to_ads_sfixed( 0.23176), im => to_ads_sfixed(-0.71329) ),
			( re => to_ads_sfixed( 0.24241), im => to_ads_sfixed(-0.70975) ),
			( re => to_ads_sfixed( 0.25300), im => to_ads_sfixed(-0.70604) ),
			( re => to_ads_sfixed( 0.26353), im => to_ads_sfixed(-0.70218) ),
			( re => to_ads_sfixed( 0.27401), im => to_ads_sfixed(-0.69816) ),
			( re => to_ads_sfixed( 0.28442), im => to_ads_sfixed(-0.69398) ),
			( re => to_ads_sfixed( 0.29477), im => to_ads_sfixed(-0.68965) ),
			( re => to_ads_sfixed( 0.30505), im => to_ads_sfixed(-0.68516) ),
			( re => to_ads_sfixed( 0.31527), im => to_ads_sfixed(-0.68052) ),
			( re => to_ads_sfixed( 0.32541), im => to_ads_sfixed(-0.67573) ),
			( re => to_ads_sfixed( 0.33548), im => to_ads_sfixed(-0.67078) ),
			( re => to_ads_sfixed( 0.34548), im => to_ads_sfixed(-0.66569) ),
			( re => to_ads_sfixed( 0.35540), im => to_ads_sfixed(-0.66045) ),
			( re => to_ads_sfixed( 0.36524), im => to_ads_sfixed(-0.65506) ),
			( re => to_ads_sfixed( 0.37500), im => to_ads_sfixed(-0.64952) ),
			( re => to_ads_sfixed( 0.38467), im => to_ads_sfixed(-0.64384) ),
			( re => to_ads_sfixed( 0.39426), im => to_ads_sfixed(-0.63801) ),
			( re => to_ads_sfixed( 0.40376), im => to_ads_sfixed(-0.63204) ),
			( re => to_ads_sfixed( 0.41317), im => to_ads_sfixed(-0.62593) ),
			( re => to_ads_sfixed( 0.42249), im => to_ads_sfixed(-0.61968) ),
			( re => to_ads_sfixed( 0.43171), im => to_ads_sfixed(-0.61329) ),
			( re => to_ads_sfixed( 0.44084), im => to_ads_sfixed(-0.60676) ),
			( re => to_ads_sfixed( 0.44987), im => to_ads_sfixed(-0.60010) ),
			( re => to_ads_sfixed( 0.45879), im => to_ads_sfixed(-0.59330) ),
			( re => to_ads_sfixed( 0.46762), im => to_ads_sfixed(-0.58637) ),
			( re => to_ads_sfixed( 0.47634), im => to_ads_sfixed(-0.57931) ),
			( re => to_ads_sfixed( 0.48495), im => to_ads_sfixed(-0.57212) ),
			( re => to_ads_sfixed( 0.49345), im => to_ads_sfixed(-0.56480) ),
			( re => to_ads_sfixed( 0.50185), im => to_ads_sfixed(-0.55736) ),
			( re => to_ads_sfixed( 0.51013), im => to_ads_sfixed(-0.54979) ),
			( re => to_ads_sfixed( 0.51830), im => to_ads_sfixed(-0.54210) ),
			( re => to_ads_sfixed( 0.52635), im => to_ads_sfixed(-0.53428) ),
			( re => to_ads_sfixed( 0.53428), im => to_ads_sfixed(-0.52635) ),
			( re => to_ads_sfixed( 0.54210), im => to_ads_sfixed(-0.51830) ),
			( re => to_ads_sfixed( 0.54979), im => to_ads_sfixed(-0.51013) ),
			( re => to_ads_sfixed( 0.55736), im => to_ads_sfixed(-0.50185) ),
			( re => to_ads_sfixed( 0.56480), im => to_ads_sfixed(-0.49345) ),
			( re => to_ads_sfixed( 0.57212), im => to_ads_sfixed(-0.48495) ),
			( re => to_ads_sfixed( 0.57931), im => to_ads_sfixed(-0.47634) ),
			( re => to_ads_sfixed( 0.58637), im => to_ads_sfixed(-0.46762) ),
			( re => to_ads_sfixed( 0.59330), im => to_ads_sfixed(-0.45879) ),
			( re => to_ads_sfixed( 0.60010), im => to_ads_sfixed(-0.44987) ),
			( re => to_ads_sfixed( 0.60676), im => to_ads_sfixed(-0.44084) ),
			( re => to_ads_sfixed( 0.61329), im => to_ads_sfixed(-0.43171) ),
			( re => to_ads_sfixed( 0.61968), im => to_ads_sfixed(-0.42249) ),
			( re => to_ads_sfixed( 0.62593), im => to_ads_sfixed(-0.41317) ),
			( re => to_ads_sfixed( 0.63204), im => to_ads_sfixed(-0.40376) ),
			( re => to_ads_sfixed( 0.63801), im => to_ads_sfixed(-0.39426) ),
			( re => to_ads_sfixed( 0.64384), im => to_ads_sfixed(-0.38467) ),
			( re => to_ads_sfixed( 0.64952), im => to_ads_sfixed(-0.37500) ),
			( re => to_ads_sfixed( 0.65506), im => to_ads_sfixed(-0.36524) ),
			( re => to_ads_sfixed( 0.66045), im => to_ads_sfixed(-0.35540) ),
			( re => to_ads_sfixed( 0.66569), im => to_ads_sfixed(-0.34548) ),
			( re => to_ads_sfixed( 0.67078), im => to_ads_sfixed(-0.33548) ),
			( re => to_ads_sfixed( 0.67573), im => to_ads_sfixed(-0.32541) ),
			( re => to_ads_sfixed( 0.68052), im => to_ads_sfixed(-0.31527) ),
			( re => to_ads_sfixed( 0.68516), im => to_ads_sfixed(-0.30505) ),
			( re => to_ads_sfixed( 0.68965), im => to_ads_sfixed(-0.29477) ),
			( re => to_ads_sfixed( 0.69398), im => to_ads_sfixed(-0.28442) ),
			( re => to_ads_sfixed( 0.69816), im => to_ads_sfixed(-0.27401) ),
			( re => to_ads_sfixed( 0.70218), im => to_ads_sfixed(-0.26353) ),
			( re => to_ads_sfixed( 0.70604), im => to_ads_sfixed(-0.25300) ),
			( re => to_ads_sfixed( 0.70975), im => to_ads_sfixed(-0.24241) ),
			( re => to_ads_sfixed( 0.71329), im => to_ads_sfixed(-0.23176) ),
			( re => to_ads_sfixed( 0.71668), im => to_ads_sfixed(-0.22107) ),
			( re => to_ads_sfixed( 0.71991), im => to_ads_sfixed(-0.21032) ),
			( re => to_ads_sfixed( 0.72297), im => to_ads_sfixed(-0.19953) ),
			( re => to_ads_sfixed( 0.72588), im => to_ads_sfixed(-0.18869) ),
			( re => to_ads_sfixed( 0.72862), im => to_ads_sfixed(-0.17781) ),
			( re => to_ads_sfixed( 0.73120), im => to_ads_sfixed(-0.16689) ),
			( re => to_ads_sfixed( 0.73361), im => to_ads_sfixed(-0.15593) ),
			( re => to_ads_sfixed( 0.73586), im => to_ads_sfixed(-0.14494) ),
			( re => to_ads_sfixed( 0.73795), im => to_ads_sfixed(-0.13392) ),
			( re => to_ads_sfixed( 0.73987), im => to_ads_sfixed(-0.12286) ),
			( re => to_ads_sfixed( 0.74162), im => to_ads_sfixed(-0.11178) ),
			( re => to_ads_sfixed( 0.74321), im => to_ads_sfixed(-0.10067) ),
			( re => to_ads_sfixed( 0.74464), im => to_ads_sfixed(-0.08955) ),
			( re => to_ads_sfixed( 0.74589), im => to_ads_sfixed(-0.07840) ),
			( re => to_ads_sfixed( 0.74698), im => to_ads_sfixed(-0.06723) ),
			( re => to_ads_sfixed( 0.74790), im => to_ads_sfixed(-0.05605) ),
			( re => to_ads_sfixed( 0.74866), im => to_ads_sfixed(-0.04485) ),
			( re => to_ads_sfixed( 0.74924), im => to_ads_sfixed(-0.03365) ),
			( re => to_ads_sfixed( 0.74966), im => to_ads_sfixed(-0.02244) ),
			( re => to_ads_sfixed( 0.74992), im => to_ads_sfixed(-0.01122) )
		);
		
	constant seed_rom_total: natural := seed_rom'length;
	subtype seed_index_type is natural range 0 to seed_rom_total - 1;
	
	function get_next_seed_index (
			index: in seed_index_type
	) return seed_index_type;
end package seed_table;

package body seed_table is
	function get_next_seed_index (
			index: in seed_index_type
	) return seed_index_type
	is
	begin
		if index = index'high then
			return 0;
		end if;
		return index + 1;
	end function get_next_seed_index;
end package body seed_table;
